`include <mux.sv>
`include <./fetch/top_fetch.sv>
`include <./decode/top_decode.sv>
`include <./execute/top_execute.sv>
`include <./memory/top_memory.sv>
`include <./memory/inst_mem.sv>


module top #(
    parameter   DATA_WIDTH = 32
) (
    input   logic clk,
    input   logic rst,
    output  logic [DATA_WIDTH-1:0] a0    
);


    logic [DATA_WIDTH-1:0]      pc;
    logic [DATA_WIDTH-1:0]      ImmExt;
    logic                       PCSrc;
    logic [DATA_WIDTH-1:0]      instr;
    logic                       branch_l;
    logic [2:0]                 ALUctrl;
    logic                       RegWrite;
    logic                       ALUSrc;
    logic                       MemWrite;
    logic                       MemRead;
    logic                       ResultSrc;
    logic [DATA_WIDTH-1:0]      ALUResult;
    logic [DATA_WIDTH-1:0]      WriteData;
    logic [DATA_WIDTH-1:0]      Result;

    top_fetch fetch(
        .clk         (clk),
        .rst         (rst),
        .PCSrc       (PCSrc),
        .ImmExt      (ImmExt),
        .pc          (pc)
    );

    inst_mem inst_mem (
        .addr       (pc),
        .dout       (instr)
    );

    top_decode decode(
        .instr      (instr),
        .branch_l   (branch_l),
        .ALUctrl    (ALUctrl),
        .RegWrite   (RegWrite),
        .ALUSrc     (ALUSrc),
        .MemWrite   (MemWrite),
        .MemRead    (MemRead),
        .ResultSrc  (ResultSrc),
        .PCSrc      (PCSrc),
        .ImmExt     (ImmExt)
    );

    top_execute execute(
        .clk        (clk),
        .instr_11_7 (instr[11:7]),
        .instr_19_15(instr[19:15]),
        .instr_24_20(instr[24:20]),
        .ALUctrl    (ALUctrl),
        .ALUSrc     (ALUSrc),
        .WE3        (RegWrite),
        .Result     (Result),
        .ImmExt     (ImmExt),
        .a0         (a0),
        .ALUResult  (ALUResult),
        .branch_l   (branch_l),
        .WriteData  (WriteData)
    );

    top_memory memory(
        .clk        (clk), 
        .ALUResult  (ALUResult),
        .WriteData  (WriteData),
        .ResultSrc  (ResultSrc),
        .MemWrite   (MemWrite),
        .MemRead    (MemRead),
        .Result     (Result),
        .funct3     (instr[14:12])
    );

    //assign a0 = 32'd5;

endmodule
