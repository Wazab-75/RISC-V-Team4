`ifndef DEF_SV
`define DEF_SV

`define ALU_OPCODE_ADD              3'b000
`define ALU_OPCODE_SUB              3'b001
`define ALU_OPCODE_AND              3'b010
`define ALU_OPCODE_OR               3'b011
`define ALU_OPCODE_SLT              3'b101

`endif
